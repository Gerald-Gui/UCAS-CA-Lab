module tlb #()();

endmodule
