module cache();

endmodule
